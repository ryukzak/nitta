// The attributes of the buffer
parameter INVALID        = 0;
parameter VALID          = 1;
parameter SPI_FINISH     = 2;
parameter FULL           = 3;