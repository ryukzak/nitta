// megafunction wizard: %LPM_DIVIDE%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DIVIDE 

// ============================================================
// File Name: div.v
// Megafunction Name(s):
// 			LPM_DIVIDE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.1.0 Build 590 10/25/2017 SJ Lite Edition
// ************************************************************


//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module div (
	clock,
	denom,
	numer,
	quotient,
	remain);

	input	  clock;
	input	 [31:0] denom;
	input	 [31:0] numer;
	output [31:0] quotient;
	output [31:0] remain;

	parameter PIPELINE = 4;
	reg [31:0] buf_quotient[PIPELINE-1:0];
	reg [31:0] buf_remain[PIPELINE-1:0];
	wire [31:0] quotient = buf_quotient[3];
	wire [31:0] remain = buf_remain[3];

	always @(posedge clock) begin
		buf_quotient[0] <= numer / denom;
		buf_quotient[1] <= buf_quotient[0];
		buf_quotient[2] <= buf_quotient[1];
		buf_quotient[3] <= buf_quotient[2];

		buf_remain[0] <= numer % denom;
		buf_remain[1] <= buf_remain[0];
		buf_remain[2] <= buf_remain[1];
		buf_remain[3] <= buf_remain[2];
	end




endmodule
